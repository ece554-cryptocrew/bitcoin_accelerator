// test bench for an accelerator

module accel_tb ();

// accelerator outputs
logic hash_done;
logic mem_acc_read_en;
logic mem_acc_write_en;
logic [15:0] mem_acc_write_addr;
logic [15:0] mem_acc_read_addr;
logic [31:0] mem_acc_write_data;
logic [255:0] hash;


// accelerator inputs
logic mem_listen_en;
logic mem_acc_write_done;
logic mem_acc_read_data_valid;
logic [15:0] mem_listen_addr;
logic [31:0] mem_listen_data;
logic [511:0] mem_acc_read_data;
logic clk, rst_n;

// file handlers
// f1: stores randomly generated block headers
// f2: stores the SHA-256 hashes (generated by the accelerator)
//     of the headers in f1
integer f1, f2;

// block header
logic [511:0] temp_0; // applied at stage 1
logic [511:0] temp_1; // applied at stage 2


accel accel0 (.hash_done(hash_done), .hash(hash), // output
              .mem_acc_read_addr(mem_acc_read_addr),
              .mem_acc_read_en(mem_acc_read_en),
              .mem_acc_write_en(mem_acc_write_en),
              .mem_acc_write_data(mem_acc_write_data),
              .mem_acc_write_addr(mem_acc_write_addr),
             
              .mem_listen_addr(mem_listen_addr), // input
              .mem_listen_en(mem_listen_en),
              .mem_listen_data(mem_listen_data),
              .mem_acc_read_data(mem_acc_read_data),
              .mem_acc_read_data_valid(mem_acc_read_data_valid),
              .mem_acc_write_done(mem_acc_write_done),
              .clk(clk), .rst_n(rst_n)
             );


// generate random block headers(raw)
class blk_hdr_t;
    rand bit [639:0] blk_hdr;
endclass

blk_hdr_t new_blk = new();


// clock
initial clk = 0;
always
    #5 clk = ~clk;


//// testing ////
initial begin
f1 = $fopen("hash_in.txt", "w");
f2 = $fopen("simu_out_accel.txt", "w");

// reset
rst_n = 0;
mem_listen_en = 0;
mem_acc_write_done = 0;
mem_acc_read_data_valid = 0;
mem_listen_addr = 0;
mem_listen_data = 0;
mem_acc_read_data = 0;

@(negedge clk);
rst_n = 1;
@(posedge clk);

for (int k = 0; k < 1000; k++) begin

    if (new_blk.randomize() == 0)
        $display("failed to generate random number\n");
    
    $fwrite(f1, "%h\n", new_blk.blk_hdr);
    $display("raw block header = %h\n", new_blk.blk_hdr);

    {temp_0, temp_1} = {new_blk.blk_hdr, 1'b1, 319'b0, 64'b10_1000_0000};
    
    ///////////////////////////////
    ////////////Stage 1////////////
    @(posedge clk); // @ IDLE
    // start hashing
    mem_listen_en = 1;
    mem_listen_addr = 16'h5000;
    mem_listen_data = 32'b1;

    @(posedge clk); #1;// @ READ_MSG_1
    mem_listen_en = 0;
    assert (mem_acc_read_en == 1) 
    else   $error("error: mem_acc_read_en");
    assert (mem_acc_read_addr == 16'h1000) 
    else   $error("error: mem_acc_read_addr");

    // simulate reading from data memory
    repeat(3) @(posedge clk); // @ READ_MSG_1
    mem_acc_read_data_valid = 1;
    mem_acc_read_data = temp_0;

    @(posedge clk); #1;// @ WR_BUSY
    mem_acc_read_data_valid = 0;
    assert (mem_acc_write_en == 1) 
    else   $error("error: mem_acc_write_en");
    assert (mem_acc_write_addr == 16'h5000) 
    else   $error("error: mem_acc_write_addr");

    // simulate writing status bits to data memory
    repeat(3) @(posedge clk); // @ WR_BUSY
    mem_acc_write_done = 1;

    @(posedge clk); // @ INIT
    mem_acc_write_done = 0;

    @(posedge clk); // @ UPD1
    @(posedge clk); // @ HASH
    repeat(64) @(posedge clk); // @ HASH
    @(posedge clk); // @ UPD2
    @(posedge clk); // @ DONE
    ////////////Stage 1////////////
    ///////////////////////////////

    ///////////////////////////////
    ////////////Stage 2////////////
    @(posedge clk); #1; // @ READ_MSG_2
    assert (mem_acc_read_en == 1) 
    else   $error("error: mem_acc_read_en");
    assert (mem_acc_read_addr == 16'h1000) 
    else   $error("error: mem_acc_read_addr");
    
    // simulate reading from data memory
    repeat(3) @(posedge clk); // @ READ_MSG_2
    mem_acc_read_data_valid = 1;
    mem_acc_read_data = temp_1;

    @(posedge clk); // @ UPD1
    mem_acc_read_data_valid = 0;
    @(posedge clk); // @ HASH
    repeat(64) @(posedge clk); // @ HASH
    @(posedge clk); // @ UPD2
    @(posedge clk); // @ DONE
    ////////////Stage 2////////////
    ///////////////////////////////

    ///////////////////////////////
    ////////////Stage 3////////////
    @(posedge clk); // @ INIT
    @(posedge clk); // @ UPD1
    @(posedge clk); // @ HASH
    repeat(64) @(posedge clk); // @ HASH
    @(posedge clk); // @ UPD2
    @(posedge clk); // @ DONE
    ////////////Stage 3////////////
    ///////////////////////////////

    ///////////////////////////////
    ///////////Write Back//////////
    @(posedge clk); #1 // @ WRITE_H0
    assert (hash_done == 1)
    else   $error("error: hash_done");
    $display("final hash = %h\n", hash);
    $fwrite(f2, "%h\n", hash);
    // simulate writing hash value to data memory
    repeat(3) @(posedge clk); // @ WRITE_H0
    // **** write_done can only be asserted for 1 cycle
    mem_acc_write_done = 1;
    @(posedge clk); // @ WRITE_H1
    mem_acc_write_done = 0;
    repeat(3) @(posedge clk); // @ WRITE_H1
    mem_acc_write_done = 1;
    @(posedge clk); // @ WRITE_H2
    mem_acc_write_done = 0;
    repeat(3) @(posedge clk); // @ WRITE_H2
    mem_acc_write_done = 1;
    @(posedge clk); // @ WRITE_H3
    mem_acc_write_done = 0;
    repeat(3) @(posedge clk); // @ WRITE_H3
    mem_acc_write_done = 1;
    @(posedge clk); // @ WRITE_H4
    mem_acc_write_done = 0;
    repeat(3) @(posedge clk); // @ WRITE_H4
    mem_acc_write_done = 1;
    @(posedge clk); // @ WRITE_H5
    mem_acc_write_done = 0;
    repeat(3) @(posedge clk); // @ WRITE_H5
    mem_acc_write_done = 1;
    @(posedge clk); // @ WRITE_H6
    mem_acc_write_done = 0;
    repeat(3) @(posedge clk); // @ WRITE_H6
    mem_acc_write_done = 1;
    @(posedge clk); // @ WRITE_H7
    mem_acc_write_done = 0;
    repeat(3) @(posedge clk); // @ WRITE_H7
    mem_acc_write_done = 1;
    @(posedge clk); // @ WR_DONE
    mem_acc_write_done = 0;
    repeat(3) @(posedge clk); // @ WR_DONE
    mem_acc_write_done = 1;
    @(posedge clk); // @ IDLE
    mem_acc_write_done = 0;
    ///////////Write Back//////////
    ///////////////////////////////
end // end for

$fclose(f1);
$fclose(f2);
$stop;

end // end initial
//// end testing ////


endmodule

