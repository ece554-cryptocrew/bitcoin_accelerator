module cpu_alu(A,B,Op,Flags,Out);

input [31:0] A;
input [31:0] B;
input [7:0] Op;
output [31:0] Flags;
output [31:0] Out;

logic [31:0] top42muxOut;
logic [31:0] bot42muxOut;
logic [31:0] bPassthrough;
logic [31:0] rotateOut; 
logic [31:0] topFinalMuxOut;
logic [31:0] bottomFinalMuxOut;


assign bPassthrough = Op[2] ? (A + B) : B; // Mux on diagram with Op[2]
assign top42muxOut = Op[2] ? (A * B) : Op[1] ? (A - B) : (A + B); // Top 4:2 mux.  If Op[2:1] is 3 or 2, then Mult, if 1, Sub, if 0 add
assign bot42muxOut = Op[2] ? rotateOut : Op[1] ? (A >> B) : (A << B); // Bot 4:2 mux.  If Op[2:1] is 3 or 2 then rotate by B etc..
assign topFinalMuxOut = Op[4] ? top42muxOut : bot42muxOut;
assign bottomFinalMuxOut = Op[7] ? (Op[2] ? (A+B) : B) : A;
assign Out = (Op[4] || Op[5]) ? topFinalMuxOut : bottomFinalMuxOut;

always_comb begin

case(B[4:0])
	5'h0: rotateOut = A;
	5'h1: rotateOut = {A[0],A[31:1]};
	5'h2: rotateOut = {A[1:0],A[31:2]};
	5'h3: rotateOut = {A[2:0],A[31:3]};
	5'h4: rotateOut = {A[3:0],A[31:4]};
	5'h5: rotateOut = {A[4:0],A[31:5]};
	5'h6: rotateOut = {A[5:0],A[31:6]};
	5'h7: rotateOut = {A[6:0],A[31:7]};
	5'h8: rotateOut = {A[7:0],A[31:8]};
	5'h9: rotateOut = {A[8:0],A[31:9]};
	5'd10: rotateOut = {A[9:0],A[31:10]};
	5'd11: rotateOut = {A[10:0],A[31:11]};
	5'd12: rotateOut = {A[11:0],A[31:12]};
	5'd13: rotateOut = {A[12:0],A[31:13]};
	5'd14: rotateOut = {A[13:0],A[31:14]};
	5'd15: rotateOut = {A[14:0],A[31:15]};
	5'd16: rotateOut = {A[15:0],A[31:16]};
	5'd17: rotateOut = {A[16:0],A[31:17]};
	5'd18: rotateOut = {A[17:0],A[31:18]};
	5'd19: rotateOut = {A[18:0],A[31:19]};
	5'd20: rotateOut = {A[19:0],A[31:20]};
	5'd21: rotateOut = {A[20:0],A[31:21]};
	5'd22: rotateOut = {A[21:0],A[31:22]};
	5'd23: rotateOut = {A[22:0],A[31:23]};
	5'd24: rotateOut = {A[23:0],A[31:24]};
	5'd25: rotateOut = {A[24:0],A[31:25]};
	5'd26: rotateOut = {A[25:0],A[31:26]};
	5'd27: rotateOut = {A[26:0],A[31:27]};
	5'd28: rotateOut = {A[27:0],A[31:28]};
	5'd29: rotateOut = {A[28:0],A[31:29]};
	5'd30: rotateOut = {A[29:0],A[31:30]};
	5'd31: rotateOut = {A[30:0],A[31]};
endcase

end

endmodule
